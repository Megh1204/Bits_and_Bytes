`timescale 1ns / 1ps

module testbench();

reg [63:0] in;
wire out;

unknown_x_detector inst(
    .in(in),
    .out(out)
    );
    
initial begin
    in = 64'b0;
    #10
    in = 64'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    //out = 0;
    #10
    in = 64'b0000_0000_0000_0x00_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    //out = x;
    #50
    in = 64'b0000_0000_0000_1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
    //out = 1;
    #50
    $stop;
end 

endmodule
